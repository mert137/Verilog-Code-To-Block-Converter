module case2_block (
input port_in_0,
input port_in_1,
output port_out_2,
output port_out_3,
inout port_inout_4
);
endmodule
